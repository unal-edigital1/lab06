`timescale 1ns / 1ps

module FSM_game (
	 	input clk,
		input rst,
		input in1,
		input in2,
		output mem_px_addr,
		output mem_px_data,
		output px_wr
   );

	/**aca va el codigo de cada grupo**/
endmodule
